library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.edc_common.all;

package interpolator_common is
    type interpolator_input_tran is record
        infr : complex10;  
        supr : complex10;  
    end record;

    type interpolator_output_tran_type is array (0 to 11) of complex10;

    type interpolator_output_tran is record
        data : interpolator_output_tran_type;
    end record;

    function interpolator_predict(
        input_tran : interpolator_input_tran
    ) return interpolator_output_tran;

end package interpolator_common;

package body interpolator_common is

    function interpolator_predict(
        input_tran : interpolator_input_tran
    ) return interpolator_output_tran is
        variable output_tran : interpolator_output_tran;
        variable infr_re, infr_im : integer;
        variable supr_re, supr_im : integer;
    begin
        infr_re := to_integer(input_tran.infr.re);
        infr_im := to_integer(input_tran.infr.im);
        supr_re := to_integer(input_tran.supr.re);
        supr_im := to_integer(input_tran.supr.im);

        for i in 0 to 11 loop
            output_tran.data(i).re :=  to_signed( (infr_re * (12 - i)/12 + supr_re * i/12) * 3/4, 10);
            output_tran.data(i).im :=  to_signed( (infr_im * (12 - i)/12 + supr_im * i/12) * 3/4, 10);
        end loop;

        return output_tran;
    end function;
    
end package body interpolator_common;
