library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.types_pkg.all;

entity sigmoid is
    port (
        x : in  q8_8;   -- Q8.8 input, between -8.0 y +8.0
        y : out q8_8    -- sigmoid(x) output in Q8.8
    );
end sigmoid;

architecture rtl of sigmoid is
    type lut_array is array(0 to 255) of q8_8;

    constant lut : lut_array := (
        to_signed(0, 16),  -- x"0000"  sig(-8.0000) = 0.000000
        to_signed(0, 16),  -- x"0000"  sig(-7.9373) = 0.000000
        to_signed(0, 16),  -- x"0000"  sig(-7.8745) = 0.000000
        to_signed(0, 16),  -- x"0000"  sig(-7.8118) = 0.000000
        to_signed(0, 16),  -- x"0000"  sig(-7.7490) = 0.000000
        to_signed(0, 16),  -- x"0000"  sig(-7.6863) = 0.000000
        to_signed(0, 16),  -- x"0000"  sig(-7.6235) = 0.000000
        to_signed(0, 16),  -- x"0000"  sig(-7.5608) = 0.000000
        to_signed(0, 16),  -- x"0000"  sig(-7.4980) = 0.000000
        to_signed(0, 16),  -- x"0000"  sig(-7.4353) = 0.000000
        to_signed(0, 16),  -- x"0000"  sig(-7.3725) = 0.000000
        to_signed(0, 16),  -- x"0000"  sig(-7.3098) = 0.000000
        to_signed(0, 16),  -- x"0000"  sig(-7.2471) = 0.000000
        to_signed(0, 16),  -- x"0000"  sig(-7.1843) = 0.000000
        to_signed(0, 16),  -- x"0000"  sig(-7.1216) = 0.000000
        to_signed(0, 16),  -- x"0000"  sig(-7.0588) = 0.000000
        to_signed(0, 16),  -- x"0000"  sig(-6.9961) = 0.000000
        to_signed(0, 16),  -- x"0000"  sig(-6.9333) = 0.000000
        to_signed(0, 16),  -- x"0000"  sig(-6.8706) = 0.000000
        to_signed(0, 16),  -- x"0000"  sig(-6.8078) = 0.000000
        to_signed(0, 16),  -- x"0000"  sig(-6.7451) = 0.000000
        to_signed(0, 16),  -- x"0000"  sig(-6.6824) = 0.000000
        to_signed(0, 16),  -- x"0000"  sig(-6.6196) = 0.000000
        to_signed(0, 16),  -- x"0000"  sig(-6.5569) = 0.000000
        to_signed(0, 16),  -- x"0000"  sig(-6.4941) = 0.000000
        to_signed(0, 16),  -- x"0000"  sig(-6.4314) = 0.000000
        to_signed(0, 16),  -- x"0000"  sig(-6.3686) = 0.000000
        to_signed(0, 16),  -- x"0000"  sig(-6.3059) = 0.000000
        to_signed(0, 16),  -- x"0000"  sig(-6.2431) = 0.000000
        to_signed(1, 16),  -- x"0001"  sig(-6.1804) = 0.003906
        to_signed(1, 16),  -- x"0001"  sig(-6.1176) = 0.003906
        to_signed(1, 16),  -- x"0001"  sig(-6.0549) = 0.003906
        to_signed(1, 16),  -- x"0001"  sig(-5.9922) = 0.003906
        to_signed(1, 16),  -- x"0001"  sig(-5.9294) = 0.003906
        to_signed(1, 16),  -- x"0001"  sig(-5.8667) = 0.003906
        to_signed(1, 16),  -- x"0001"  sig(-5.8039) = 0.003906
        to_signed(1, 16),  -- x"0001"  sig(-5.7412) = 0.003906
        to_signed(1, 16),  -- x"0001"  sig(-5.6784) = 0.003906
        to_signed(1, 16),  -- x"0001"  sig(-5.6157) = 0.003906
        to_signed(1, 16),  -- x"0001"  sig(-5.5529) = 0.003906
        to_signed(1, 16),  -- x"0001"  sig(-5.4902) = 0.003906
        to_signed(1, 16),  -- x"0001"  sig(-5.4275) = 0.003906
        to_signed(1, 16),  -- x"0001"  sig(-5.3647) = 0.003906
        to_signed(1, 16),  -- x"0001"  sig(-5.3020) = 0.003906
        to_signed(1, 16),  -- x"0001"  sig(-5.2392) = 0.003906
        to_signed(1, 16),  -- x"0001"  sig(-5.1765) = 0.003906
        to_signed(2, 16),  -- x"0002"  sig(-5.1137) = 0.007812
        to_signed(2, 16),  -- x"0002"  sig(-5.0510) = 0.007812
        to_signed(2, 16),  -- x"0002"  sig(-4.9882) = 0.007812
        to_signed(2, 16),  -- x"0002"  sig(-4.9255) = 0.007812
        to_signed(2, 16),  -- x"0002"  sig(-4.8627) = 0.007812
        to_signed(2, 16),  -- x"0002"  sig(-4.8000) = 0.007812
        to_signed(2, 16),  -- x"0002"  sig(-4.7373) = 0.007812
        to_signed(2, 16),  -- x"0002"  sig(-4.6745) = 0.007812
        to_signed(3, 16),  -- x"0003"  sig(-4.6118) = 0.011719
        to_signed(3, 16),  -- x"0003"  sig(-4.5490) = 0.011719
        to_signed(3, 16),  -- x"0003"  sig(-4.4863) = 0.011719
        to_signed(3, 16),  -- x"0003"  sig(-4.4235) = 0.011719
        to_signed(3, 16),  -- x"0003"  sig(-4.3608) = 0.011719
        to_signed(3, 16),  -- x"0003"  sig(-4.2980) = 0.011719
        to_signed(4, 16),  -- x"0004"  sig(-4.2353) = 0.015625
        to_signed(4, 16),  -- x"0004"  sig(-4.1725) = 0.015625
        to_signed(4, 16),  -- x"0004"  sig(-4.1098) = 0.015625
        to_signed(4, 16),  -- x"0004"  sig(-4.0471) = 0.015625
        to_signed(5, 16),  -- x"0005"  sig(-3.9843) = 0.019531
        to_signed(5, 16),  -- x"0005"  sig(-3.9216) = 0.019531
        to_signed(5, 16),  -- x"0005"  sig(-3.8588) = 0.019531
        to_signed(6, 16),  -- x"0006"  sig(-3.7961) = 0.023438
        to_signed(6, 16),  -- x"0006"  sig(-3.7333) = 0.023438
        to_signed(6, 16),  -- x"0006"  sig(-3.6706) = 0.023438
        to_signed(7, 16),  -- x"0007"  sig(-3.6078) = 0.027344
        to_signed(7, 16),  -- x"0007"  sig(-3.5451) = 0.027344
        to_signed(8, 16),  -- x"0008"  sig(-3.4824) = 0.031250
        to_signed(8, 16),  -- x"0008"  sig(-3.4196) = 0.031250
        to_signed(9, 16),  -- x"0009"  sig(-3.3569) = 0.035156
        to_signed(9, 16),  -- x"0009"  sig(-3.2941) = 0.035156
        to_signed(10, 16),  -- x"000A"  sig(-3.2314) = 0.039062
        to_signed(10, 16),  -- x"000A"  sig(-3.1686) = 0.039062
        to_signed(11, 16),  -- x"000B"  sig(-3.1059) = 0.042969
        to_signed(12, 16),  -- x"000C"  sig(-3.0431) = 0.046875
        to_signed(12, 16),  -- x"000C"  sig(-2.9804) = 0.046875
        to_signed(13, 16),  -- x"000D"  sig(-2.9176) = 0.050781
        to_signed(14, 16),  -- x"000E"  sig(-2.8549) = 0.054688
        to_signed(15, 16),  -- x"000F"  sig(-2.7922) = 0.058594
        to_signed(16, 16),  -- x"0010"  sig(-2.7294) = 0.062500
        to_signed(17, 16),  -- x"0011"  sig(-2.6667) = 0.066406
        to_signed(18, 16),  -- x"0012"  sig(-2.6039) = 0.070312
        to_signed(19, 16),  -- x"0013"  sig(-2.5412) = 0.074219
        to_signed(20, 16),  -- x"0014"  sig(-2.4784) = 0.078125
        to_signed(21, 16),  -- x"0015"  sig(-2.4157) = 0.082031
        to_signed(22, 16),  -- x"0016"  sig(-2.3529) = 0.085938
        to_signed(24, 16),  -- x"0018"  sig(-2.2902) = 0.093750
        to_signed(25, 16),  -- x"0019"  sig(-2.2275) = 0.097656
        to_signed(26, 16),  -- x"001A"  sig(-2.1647) = 0.101562
        to_signed(28, 16),  -- x"001C"  sig(-2.1020) = 0.109375
        to_signed(29, 16),  -- x"001D"  sig(-2.0392) = 0.113281
        to_signed(31, 16),  -- x"001F"  sig(-1.9765) = 0.121094
        to_signed(33, 16),  -- x"0021"  sig(-1.9137) = 0.128906
        to_signed(35, 16),  -- x"0023"  sig(-1.8510) = 0.136719
        to_signed(37, 16),  -- x"0025"  sig(-1.7882) = 0.144531
        to_signed(39, 16),  -- x"0027"  sig(-1.7255) = 0.152344
        to_signed(41, 16),  -- x"0029"  sig(-1.6627) = 0.160156
        to_signed(43, 16),  -- x"002B"  sig(-1.6000) = 0.167969
        to_signed(45, 16),  -- x"002D"  sig(-1.5373) = 0.175781
        to_signed(48, 16),  -- x"0030"  sig(-1.4745) = 0.187500
        to_signed(50, 16),  -- x"0032"  sig(-1.4118) = 0.195312
        to_signed(53, 16),  -- x"0035"  sig(-1.3490) = 0.207031
        to_signed(55, 16),  -- x"0037"  sig(-1.2863) = 0.214844
        to_signed(58, 16),  -- x"003A"  sig(-1.2235) = 0.226562
        to_signed(61, 16),  -- x"003D"  sig(-1.1608) = 0.238281
        to_signed(64, 16),  -- x"0040"  sig(-1.0980) = 0.250000
        to_signed(67, 16),  -- x"0043"  sig(-1.0353) = 0.261719
        to_signed(70, 16),  -- x"0046"  sig(-0.9725) = 0.273438
        to_signed(73, 16),  -- x"0049"  sig(-0.9098) = 0.285156
        to_signed(77, 16),  -- x"004D"  sig(-0.8471) = 0.300781
        to_signed(80, 16),  -- x"0050"  sig(-0.7843) = 0.312500
        to_signed(84, 16),  -- x"0054"  sig(-0.7216) = 0.328125
        to_signed(87, 16),  -- x"0057"  sig(-0.6588) = 0.339844
        to_signed(91, 16),  -- x"005B"  sig(-0.5961) = 0.355469
        to_signed(95, 16),  -- x"005F"  sig(-0.5333) = 0.371094
        to_signed(98, 16),  -- x"0062"  sig(-0.4706) = 0.382812
        to_signed(102, 16),  -- x"0066"  sig(-0.4078) = 0.398438
        to_signed(106, 16),  -- x"006A"  sig(-0.3451) = 0.414062
        to_signed(110, 16),  -- x"006E"  sig(-0.2824) = 0.429688
        to_signed(114, 16),  -- x"0072"  sig(-0.2196) = 0.445312
        to_signed(118, 16),  -- x"0076"  sig(-0.1569) = 0.460938
        to_signed(122, 16),  -- x"007A"  sig(-0.0941) = 0.476562
        to_signed(126, 16),  -- x"007E"  sig(-0.0314) = 0.492188
        to_signed(130, 16),  -- x"0082"  sig(0.0314) = 0.507812
        to_signed(134, 16),  -- x"0086"  sig(0.0941) = 0.523438
        to_signed(138, 16),  -- x"008A"  sig(0.1569) = 0.539062
        to_signed(142, 16),  -- x"008E"  sig(0.2196) = 0.554688
        to_signed(146, 16),  -- x"0092"  sig(0.2824) = 0.570312
        to_signed(150, 16),  -- x"0096"  sig(0.3451) = 0.585938
        to_signed(154, 16),  -- x"009A"  sig(0.4078) = 0.601562
        to_signed(158, 16),  -- x"009E"  sig(0.4706) = 0.617188
        to_signed(161, 16),  -- x"00A1"  sig(0.5333) = 0.628906
        to_signed(165, 16),  -- x"00A5"  sig(0.5961) = 0.644531
        to_signed(169, 16),  -- x"00A9"  sig(0.6588) = 0.660156
        to_signed(172, 16),  -- x"00AC"  sig(0.7216) = 0.671875
        to_signed(176, 16),  -- x"00B0"  sig(0.7843) = 0.687500
        to_signed(179, 16),  -- x"00B3"  sig(0.8471) = 0.699219
        to_signed(183, 16),  -- x"00B7"  sig(0.9098) = 0.714844
        to_signed(186, 16),  -- x"00BA"  sig(0.9725) = 0.726562
        to_signed(189, 16),  -- x"00BD"  sig(1.0353) = 0.738281
        to_signed(192, 16),  -- x"00C0"  sig(1.0980) = 0.750000
        to_signed(195, 16),  -- x"00C3"  sig(1.1608) = 0.761719
        to_signed(198, 16),  -- x"00C6"  sig(1.2235) = 0.773438
        to_signed(201, 16),  -- x"00C9"  sig(1.2863) = 0.785156
        to_signed(203, 16),  -- x"00CB"  sig(1.3490) = 0.792969
        to_signed(206, 16),  -- x"00CE"  sig(1.4118) = 0.804688
        to_signed(208, 16),  -- x"00D0"  sig(1.4745) = 0.812500
        to_signed(211, 16),  -- x"00D3"  sig(1.5373) = 0.824219
        to_signed(213, 16),  -- x"00D5"  sig(1.6000) = 0.832031
        to_signed(215, 16),  -- x"00D7"  sig(1.6627) = 0.839844
        to_signed(217, 16),  -- x"00D9"  sig(1.7255) = 0.847656
        to_signed(219, 16),  -- x"00DB"  sig(1.7882) = 0.855469
        to_signed(221, 16),  -- x"00DD"  sig(1.8510) = 0.863281
        to_signed(223, 16),  -- x"00DF"  sig(1.9137) = 0.871094
        to_signed(225, 16),  -- x"00E1"  sig(1.9765) = 0.878906
        to_signed(227, 16),  -- x"00E3"  sig(2.0392) = 0.886719
        to_signed(228, 16),  -- x"00E4"  sig(2.1020) = 0.890625
        to_signed(230, 16),  -- x"00E6"  sig(2.1647) = 0.898438
        to_signed(231, 16),  -- x"00E7"  sig(2.2275) = 0.902344
        to_signed(232, 16),  -- x"00E8"  sig(2.2902) = 0.906250
        to_signed(234, 16),  -- x"00EA"  sig(2.3529) = 0.914062
        to_signed(235, 16),  -- x"00EB"  sig(2.4157) = 0.917969
        to_signed(236, 16),  -- x"00EC"  sig(2.4784) = 0.921875
        to_signed(237, 16),  -- x"00ED"  sig(2.5412) = 0.925781
        to_signed(238, 16),  -- x"00EE"  sig(2.6039) = 0.929688
        to_signed(239, 16),  -- x"00EF"  sig(2.6667) = 0.933594
        to_signed(240, 16),  -- x"00F0"  sig(2.7294) = 0.937500
        to_signed(241, 16),  -- x"00F1"  sig(2.7922) = 0.941406
        to_signed(242, 16),  -- x"00F2"  sig(2.8549) = 0.945312
        to_signed(243, 16),  -- x"00F3"  sig(2.9176) = 0.949219
        to_signed(244, 16),  -- x"00F4"  sig(2.9804) = 0.953125
        to_signed(244, 16),  -- x"00F4"  sig(3.0431) = 0.953125
        to_signed(245, 16),  -- x"00F5"  sig(3.1059) = 0.957031
        to_signed(246, 16),  -- x"00F6"  sig(3.1686) = 0.960938
        to_signed(246, 16),  -- x"00F6"  sig(3.2314) = 0.960938
        to_signed(247, 16),  -- x"00F7"  sig(3.2941) = 0.964844
        to_signed(247, 16),  -- x"00F7"  sig(3.3569) = 0.964844
        to_signed(248, 16),  -- x"00F8"  sig(3.4196) = 0.968750
        to_signed(248, 16),  -- x"00F8"  sig(3.4824) = 0.968750
        to_signed(249, 16),  -- x"00F9"  sig(3.5451) = 0.972656
        to_signed(249, 16),  -- x"00F9"  sig(3.6078) = 0.972656
        to_signed(250, 16),  -- x"00FA"  sig(3.6706) = 0.976562
        to_signed(250, 16),  -- x"00FA"  sig(3.7333) = 0.976562
        to_signed(250, 16),  -- x"00FA"  sig(3.7961) = 0.976562
        to_signed(251, 16),  -- x"00FB"  sig(3.8588) = 0.980469
        to_signed(251, 16),  -- x"00FB"  sig(3.9216) = 0.980469
        to_signed(251, 16),  -- x"00FB"  sig(3.9843) = 0.980469
        to_signed(252, 16),  -- x"00FC"  sig(4.0471) = 0.984375
        to_signed(252, 16),  -- x"00FC"  sig(4.1098) = 0.984375
        to_signed(252, 16),  -- x"00FC"  sig(4.1725) = 0.984375
        to_signed(252, 16),  -- x"00FC"  sig(4.2353) = 0.984375
        to_signed(253, 16),  -- x"00FD"  sig(4.2980) = 0.988281
        to_signed(253, 16),  -- x"00FD"  sig(4.3608) = 0.988281
        to_signed(253, 16),  -- x"00FD"  sig(4.4235) = 0.988281
        to_signed(253, 16),  -- x"00FD"  sig(4.4863) = 0.988281
        to_signed(253, 16),  -- x"00FD"  sig(4.5490) = 0.988281
        to_signed(253, 16),  -- x"00FD"  sig(4.6118) = 0.988281
        to_signed(254, 16),  -- x"00FE"  sig(4.6745) = 0.992188
        to_signed(254, 16),  -- x"00FE"  sig(4.7373) = 0.992188
        to_signed(254, 16),  -- x"00FE"  sig(4.8000) = 0.992188
        to_signed(254, 16),  -- x"00FE"  sig(4.8627) = 0.992188
        to_signed(254, 16),  -- x"00FE"  sig(4.9255) = 0.992188
        to_signed(254, 16),  -- x"00FE"  sig(4.9882) = 0.992188
        to_signed(254, 16),  -- x"00FE"  sig(5.0510) = 0.992188
        to_signed(254, 16),  -- x"00FE"  sig(5.1137) = 0.992188
        to_signed(255, 16),  -- x"00FF"  sig(5.1765) = 0.996094
        to_signed(255, 16),  -- x"00FF"  sig(5.2392) = 0.996094
        to_signed(255, 16),  -- x"00FF"  sig(5.3020) = 0.996094
        to_signed(255, 16),  -- x"00FF"  sig(5.3647) = 0.996094
        to_signed(255, 16),  -- x"00FF"  sig(5.4275) = 0.996094
        to_signed(255, 16),  -- x"00FF"  sig(5.4902) = 0.996094
        to_signed(255, 16),  -- x"00FF"  sig(5.5529) = 0.996094
        to_signed(255, 16),  -- x"00FF"  sig(5.6157) = 0.996094
        to_signed(255, 16),  -- x"00FF"  sig(5.6784) = 0.996094
        to_signed(255, 16),  -- x"00FF"  sig(5.7412) = 0.996094
        to_signed(255, 16),  -- x"00FF"  sig(5.8039) = 0.996094
        to_signed(255, 16),  -- x"00FF"  sig(5.8667) = 0.996094
        to_signed(255, 16),  -- x"00FF"  sig(5.9294) = 0.996094
        to_signed(255, 16),  -- x"00FF"  sig(5.9922) = 0.996094
        to_signed(255, 16),  -- x"00FF"  sig(6.0549) = 0.996094
        to_signed(255, 16),  -- x"00FF"  sig(6.1176) = 0.996094
        to_signed(255, 16),  -- x"00FF"  sig(6.1804) = 0.996094
        to_signed(256, 16),  -- x"0100"  sig(6.2431) = 1.000000
        to_signed(256, 16),  -- x"0100"  sig(6.3059) = 1.000000
        to_signed(256, 16),  -- x"0100"  sig(6.3686) = 1.000000
        to_signed(256, 16),  -- x"0100"  sig(6.4314) = 1.000000
        to_signed(256, 16),  -- x"0100"  sig(6.4941) = 1.000000
        to_signed(256, 16),  -- x"0100"  sig(6.5569) = 1.000000
        to_signed(256, 16),  -- x"0100"  sig(6.6196) = 1.000000
        to_signed(256, 16),  -- x"0100"  sig(6.6824) = 1.000000
        to_signed(256, 16),  -- x"0100"  sig(6.7451) = 1.000000
        to_signed(256, 16),  -- x"0100"  sig(6.8078) = 1.000000
        to_signed(256, 16),  -- x"0100"  sig(6.8706) = 1.000000
        to_signed(256, 16),  -- x"0100"  sig(6.9333) = 1.000000
        to_signed(256, 16),  -- x"0100"  sig(6.9961) = 1.000000
        to_signed(256, 16),  -- x"0100"  sig(7.0588) = 1.000000
        to_signed(256, 16),  -- x"0100"  sig(7.1216) = 1.000000
        to_signed(256, 16),  -- x"0100"  sig(7.1843) = 1.000000
        to_signed(256, 16),  -- x"0100"  sig(7.2471) = 1.000000
        to_signed(256, 16),  -- x"0100"  sig(7.3098) = 1.000000
        to_signed(256, 16),  -- x"0100"  sig(7.3725) = 1.000000
        to_signed(256, 16),  -- x"0100"  sig(7.4353) = 1.000000
        to_signed(256, 16),  -- x"0100"  sig(7.4980) = 1.000000
        to_signed(256, 16),  -- x"0100"  sig(7.5608) = 1.000000
        to_signed(256, 16),  -- x"0100"  sig(7.6235) = 1.000000
        to_signed(256, 16),  -- x"0100"  sig(7.6863) = 1.000000
        to_signed(256, 16),  -- x"0100"  sig(7.7490) = 1.000000
        to_signed(256, 16),  -- x"0100"  sig(7.8118) = 1.000000
        to_signed(256, 16),  -- x"0100"  sig(7.8745) = 1.000000
        to_signed(256, 16),  -- x"0100"  sig(7.9373) = 1.000000
        to_signed(256, 16)  -- x"0100"  sig(8.0000) = 1.000000
    );

begin
    process(x)
        variable x_clip : integer;
        variable idx    : integer;
    begin
        if x < to_signed(-2048,16) then
            x_clip := -2048;
        elsif x > to_signed(2047,16) then
            x_clip := 2047;
        else
            x_clip := to_integer(x);
        end if;

        idx := (x_clip + 2048) / 16;

        if idx < 0 then
            idx := 0;
        elsif idx > 255 then
            idx := 255;
        end if;

        y <= lut(idx);
    end process;
end rtl;
