package minicalc_datatypes is

  type op_type is (sum, sub, mul);

end minicalc_datatypes;
